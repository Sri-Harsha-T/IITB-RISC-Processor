-- implementing bootloading logic for data path
library ieee;
library work;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.basic.all;

entity data_bootload is
	port(
		clk, reset, RX: in std_logic;
		T: in std_logic_vector(6 downto 0);
		S: out std_logic_vector(2 downto 0);
		address,data: out std_logic_vector(15 downto 0);
		enable: out std_logic
	);
end entity;

architecture data_bootload_arch of data_bootload is
	component uart_receive is 
		port(
			data: out std_logic_vector(7 downto 0); 
			received: out std_logic;
			clock,RX: in std_logic
		);
	end component;
	signal a_in, d_in, d_out, a_out: std_logic_vector(15 downto 0);
	signal uart_data, c_in, c_out: std_logic_vector(7 downto 0);
	signal a_ena, d_ena, c_ena: std_logic;
begin
	a_in <= (uart_data & "00000000") when (T(0) = '1' and T(1) = '0') 
		else std_logic_vector(unsigned(a_out) + to_unsigned(1,16)) when (T(0) = '1' and T(1) = '1')
		else std_logic_vector(unsigned(a_out(15 downto 8) & uart_data) - to_unsigned(1,16));
	a_ena <= T(0) or T(1);
	addr: my_reg
		generic map(16)
		port map(
			Din => a_in, Dout => a_out, clk => clk, ena => a_ena, clr => reset);
	
	d_in <= (uart_data & "00000000") when (T(2) = '1') 
		else (d_out(15 downto 8) & uart_data);
	d_ena <= T(3);
	dat: my_reg
		generic map(16)
		port map(
			Din => d_in, Dout => d_out, clk => clk, ena => d_ena, clr => reset);
	
	c_in <= uart_data when (T(4) = '1') else 
		std_logic_vector(unsigned(c_out) - to_unsigned(1,8));
	c_ena <= T(5);
	count: my_reg
		generic map(8)
		port map(
			Din => c_in, Dout => c_out, clk => clk, ena => c_ena, clr => reset);
	
	address <= a_out;
	data <= d_out;
	
	ena: process(clk)
	begin
		if(clk'event and clk = '1') then
			enable <= T(6);
		end if;
	end process;
	
	S(1) <= '1' when (uart_data = "00000000") else '0';
	S(2) <= '1' when (c_out = "00000000") else '0';	
	reception: uart_receive
		port map(RX => RX, clock => clk, received => S(0), data => uart_data);
			
end architecture;